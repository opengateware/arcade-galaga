mb88xx_inst : entity work.mb88xx
  port map (
    clock       => clock,
    ena         => ena,
    reset_n     => reset_n,
    r0_port_in  => r0_port_in,
    r1_port_in  => r1_port_in,
    r2_port_in  => r2_port_in,
    r3_port_in  => r3_port_in,
    r0_port_out => r0_port_out,
    r1_port_out => r1_port_out,
    r2_port_out => r2_port_out,
    r3_port_out => r3_port_out,
    k_port_in   => k_port_in,
    ol_port_out => ol_port_out,
    oh_port_out => oh_port_out,
    p_port_out  => p_port_out,
    stby_n      => stby_n,
    tc_n        => tc_n,
    irq_n       => irq_n,
    sc_in_n     => sc_in_n,
    si_n        => si_n,
    sc_out_n    => sc_out_n,
    so_n        => so_n,
    to_n        => to_n,
    rom_addr    => rom_addr,
    rom_data    => rom_data
  );
